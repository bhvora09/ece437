`ifndef FORWARDING_UNIT_IF_VH
`define FORWARDING_UNIT_IF_VH

// all types
`include "cpu_types_pkg.vh"

interface forwarding_unit_if;
    // import types
    import cpu_types_pkg::*;

    //in
    logic 


    //out
    logic



    
    modport fu (
        input 
        output 
    );

    modport tb (
        input 
        output 
    );
endinterface

`endif //FORWARDING_UNIT_IF_VH