`include "forwarding_unit_if.vh"
`include "cpu_types_pkg.vh"

module forwarding_unit_if
(
    input CLK, nRST,
    forwarding_unit_if.fu fuif
);

    import cpu_types_pkg::*;

    always_comb begin : LOG
        
    end
endmodule